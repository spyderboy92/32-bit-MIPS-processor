module inst_mem(clock,instruction,pc,inst)
input clock;
input [31:0]pc;
output [31:0] inst;
reg [31:0] instmem[31:0];
initial begin
	instmem[0]=32'b00000000000000000000000000000000;
	instmem[1]=32'b00000000000000000000000000000000;
	instmem[2]=32'b00000000000000000000000000000000;
	instmem[3]=32'b00000000000000000000000000000000;
	instmem[4]=32'b00000000000000000000000000000000;
	instmem[5]=32'b00000000000000000000000000000000;
	instmem[6]=32'b00000000000000000000000000000000;
	instmem[7]=32'b00000000000000000000000000000000;
	instmem[8]=32'b00000000000000000000000000000000;
	instmem[9]=32'b00000000000000000000000000000000;
	instmem[10]=32'b00000000000000000000000000000000;
	instmem[11]=32'b00000000000000000000000000000000;
	instmem[12]=32'b00000000000000000000000000000000;
	instmem[13]=32'b00000000000000000000000000000000;
	instmem[14]=32'b00000000000000000000000000000000;
	instmem[15]=32'b00000000000000000000000000000000;
	instmem[16]=32'b00000000000000000000000000000000;
	instmem[17]=32'b00000000000000000000000000000000;
	instmem[18]=32'b00000000000000000000000000000000;
	instmem[19]=32'b00000000000000000000000000000000;
	instmem[20]=32'b00000000000000000000000000000000;
	instmem[21]=32'b00000000000000000000000000000000;
	instmem[22]=32'b00000000000000000000000000000000;
	instmem[23]=32'b00000000000000000000000000000000;
	instmem[24]=32'b00000000000000000000000000000000;
	instmem[25]=32'b00000000000000000000000000000000;
	instmem[26]=32'b00000000000000000000000000000000;
	instmem[27]=32'b00000000000000000000000000000000;
	instmem[28]=32'b00000000000000000000000000000000;
	instmem[29]=32'b00000000000000000000000000000000;
	instmem[30]=32'b00000000000000000000000000000000;
	instmem[31]=32'b00000000000000000000000000000000;
end

always @(posedge clock)
	begin
		inst=instmem[pc];
	end
endmodule
