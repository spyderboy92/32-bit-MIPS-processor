module data_mem(clock, opcode,rt,address,out)
input [5:0]opcode;
input [31:0]address
input [31:0] rt;
input clock;
output [31:0] out;

reg [31:0] datamem[31:0];

initial begin 

	      datamem[0] = 32'b00000000000000000000000000000000;
        datamem[1] = 32'b00000000000000000000000000000000;
        datamem[2] = 32'b00000000000000000000000000000000;
        datamem[3] = 32'b00000000000000000000000000000000;
        datamem[4] = 32'b00000000000000000000000000000000;
        datamem[5] = 32'b00000000000000000000000000000000;
        datamem[6] = 32'b00000000000000000000000000000000;
        datamem[7] = 32'b00000000000000000000000000000000;
        datamem[8] = 32'b00000000000000000000000000000000;
        datamem[9] = 32'b00000000000000000000000000000000;
        datamem[10] = 32'b00000000000000000000000000000000;
        
	      datamem[11] = 32'b00000000000000000000000000000000;
        datamem[12] = 32'b00000000000000000000000000000000;
        datamem[13] = 32'b00000000000000000000000000000000;
        datamem[14] = 32'b00000000000000000000000000000000;
        datamem[15] = 32'b00000000000000000000000000000000;
        datamem[16] = 32'b00000000000000000000000000000000;
        datamem[17] = 32'b00000000000000000000000000000000;
        datamem[18] = 32'b00000000000000000000000000000000;
        datamem[19] = 32'b00000000000000000000000000000000;
	      datamem[20] = 32'b00000000000000000000000000000000;

        datamem[21] = 32'b00000000000000000000000000000000;
	      datamem[22] = 32'b00000000000000000000000000000000;
        datamem[23] = 32'b00000000000000000000000000000000;
	      datamem[24] = 32'b00000000000000000000000000000000;
        datamem[25] = 32'b00000000000000000000000000000000;
	      datamem[26] = 32'b00000000000000000000000000000000;
        datamem[27] = 32'b00000000000000000000000000000000;
	      datamem[28] = 32'b00000000000000000000000000000000;
        datamem[29] = 32'b00000000000000000000000000000000;
	      datamem[30] = 32'b00000000000000000000000000000000;
        datamem[31] = 32'b00000000000000000000000000000000;
	      datamem[32] = 32'b00000000000000000000000000000000;
end

assign out=datamem[address];
always @(posedge clock)
begin
	if(opcode==6'b101011)
	begin
	datamem[address]=out;
	end
end
always @(negedge clock)
begin
	if(opcode==6'b100011)
	begin
	rt=datamem[address];
	end
end

endmodule
